*******************************************************************
* Filename: Prelab2.cir
* Author: Mitchell Larson <larsonma@msoe.edu>
* Date: May 8, 2018
* Provides:
*	- Signal conditioning circiut that ranges a [0:400]mV signal to
*	- a [0:4000]mV signal using an LM741 opamp while providing
*  	- high pass filtering with a cut-off freqency of 2kHz and
*	- input buffering
*******************************************************************

*** Including the opamp library ***

.lib "opamp.lib"

*** Circuit Description ***
*** Simulation technique: time domain at 1K [0:400]mV ***

*** Power Supplies ***
VCC+ 1 0 DC 5.0
VCC- 2 0 DC -5.0

*** Input voltage ***
VS 3 0 AC 1.0 0.0

*** Resistors ***
R1 6 0 2K
R2 7 6 18K
Rf 5 0 8.1K

*** op-amps ***
X1 3 4 1 2 4 LM741
X2 5 6 1 2 7 LM741

*** capacitors ***
C1 4 5 10n

*** commands to spice ***
*** simulate two periods ***

.AC LIN 100 1 100K
.PROBE

.End
